library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity adder_16b is
  port ( src_a : in std_logic_vector(15 downto 0);
        src_b : in std_logic_vector(15 downto 0);
        sum : out std_logic_vector(15 downto 0);
        carry_out : out std_logic );
end adder_16b;
architecture behavioural of adder_16b is
signal sig_result : std_logic_vector(16 downto 0);
begin
  sig_result <= ('0' & src_a) + ('0' & src_b);
  sum <= sig_result(15 downto 0);
  carry_out <= sig_result(16);
end behavioural;
