----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:03:46 10/08/2017 
-- Design Name: 
-- Module Name:    nBitCounter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity nBitCounter is

	 generic(n: natural :=10);
    Port ( clk : in  STD_LOGIC;
           en : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           counterOut : out  STD_LOGIC_VECTOR(n-1 downto 0));
end nBitCounter;

architecture Behavioral of nBitCounter is

	signal counterValue: std_logic_vector(n-1 downto 0);

begin

	process(clk, en, rst)
	begin
		if rst = '1' then
			counterValue <= (others => '0');
		elsif rising_edge(clk) then
			if en = '1' then
				counterValue <= counterValue+1;
			end if;
		end if;
	end process;
	
	counterOut <= counterValue;

end Behavioral;

